`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:14:45 10/12/2016 
// Design Name: 
// Module Name:    top 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module top(
    );

bcd instance_name (
    .life(life), 
    .fenshu(fenshu), 
    .fenshu2(fenshu2), 
    .fenshu1(fenshu1), 
    .fenshu0(fenshu0), 
    .shengming(shengming)
    );

endmodule
